`define UART_MASTER_SYSCLK 5e+07
`define UART_BAUD_RATE 57600
`define LUT_BASED
