//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Sun Feb  9 17:07:40 2025

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire [23:0] prom_inst_1_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h91919191919191919191919191919191919191919191919191919191916678A1;
defparam prom_inst_0.INIT_RAM_01 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_02 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_03 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_04 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_05 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_06 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_07 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_08 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_09 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_0A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_0B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_0C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_0D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_0E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_0F = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_10 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_11 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_12 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_13 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_14 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_15 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_16 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_17 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_18 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_19 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_1A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_1B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_1C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_1D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_1E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_1F = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_20 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_21 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_22 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_23 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_24 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_25 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_26 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_27 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_28 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_29 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_2A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_2B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_2C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_2D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_2E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_2F = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_30 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_31 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_32 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_33 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_34 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_35 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_36 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_37 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_38 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_39 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_3A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_3B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_3C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_3D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_3E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_0.INIT_RAM_3F = 256'h9191919191919191919191919191919191919191919191919191919191919191;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "ASYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_08 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_09 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_0A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_0B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_0C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_0D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_0E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_0F = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_10 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_11 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_12 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_13 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_14 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_15 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_16 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_17 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_18 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_19 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_1A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_1B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_1C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_1D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_1E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_1F = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_20 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_21 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_22 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_23 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_24 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_25 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_26 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_27 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_28 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_29 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_2A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_2B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_2C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_2D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_2E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_2F = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_30 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_31 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_32 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_33 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_34 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_35 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_36 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_37 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_38 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_39 = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_3A = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_3B = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_3C = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_3D = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_3E = 256'h9191919191919191919191919191919191919191919191919191919191919191;
defparam prom_inst_1.INIT_RAM_3F = 256'h9191919191919191919191919191919191919191919191919191919191919191;

endmodule //Gowin_pROM
